module Quantizer #(
    parameter num_bit
) (
    input  [num_bit - 1:0] in,
    output [num_bit - 1:0] out
);



endmodule
